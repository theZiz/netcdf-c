netcdf input {
dimensions:
	initial_time0_hours = UNLIMITED ; // (1 currently)
	lat_0 = 205 ;
	lon_0 = 253 ;
	ncl_strlen_0 = 18 ;
variables:
	float TMP_P0_L103_GLL0(initial_time0_hours, lat_0, lon_0) ;
		TMP_P0_L103_GLL0:forecast_time_units = "hours" ;
		TMP_P0_L103_GLL0:forecast_time = 0 ;
		TMP_P0_L103_GLL0:level = 2.f ;
		TMP_P0_L103_GLL0:level_type = "Specified height level above ground (m)" ;
		TMP_P0_L103_GLL0:parameter_template_discipline_category_number = 0, 0, 0, 0 ;
		TMP_P0_L103_GLL0:parameter_discipline_and_category = "Meteorological products, Temperature" ;
		TMP_P0_L103_GLL0:grid_type = "Latitude/longitude" ;
		TMP_P0_L103_GLL0:_FillValue = 1.e+20f ;
		TMP_P0_L103_GLL0:units = "K" ;
		TMP_P0_L103_GLL0:long_name = "Temperature" ;
		TMP_P0_L103_GLL0:production_status = "Operational products" ;
		TMP_P0_L103_GLL0:center = "US National Weather Service - NCEP (WMC)" ;
	char initial_time0(initial_time0_hours, ncl_strlen_0) ;
		initial_time0:NCL_converted_from_type = "string" ;
		initial_time0:units = "mm/dd/yyyy (hh:mm)" ;
		initial_time0:long_name = "Initial time of first record" ;
	double initial_time0_encoded(initial_time0_hours) ;
		initial_time0_encoded:units = "yyyymmddhh.hh_frac" ;
		initial_time0_encoded:long_name = "initial time encoded as double" ;
	double initial_time0_hours(initial_time0_hours) ;
		initial_time0_hours:units = "hours since 1800-01-01 00:00" ;
		initial_time0_hours:long_name = "initial time" ;
	float lat_0(lat_0) ;
		lat_0:La1 = 90.f ;
		lat_0:Lo1 = 0.f ;
		lat_0:La2 = -90.f ;
		lat_0:Lo2 = 359.75f ;
		lat_0:Di = 0.25f ;
		lat_0:Dj = 0.25f ;
		lat_0:units = "degrees_north" ;
		lat_0:grid_type = "Latitude/Longitude" ;
		lat_0:long_name = "latitude" ;
	float lon_0(lon_0) ;
		lon_0:La1 = 90.f ;
		lon_0:Lo1 = 0.f ;
		lon_0:La2 = -90.f ;
		lon_0:Lo2 = 359.75f ;
		lon_0:Di = 0.25f ;
		lon_0:Dj = 0.25f ;
		lon_0:units = "degrees_east" ;
		lon_0:grid_type = "Latitude/Longitude" ;
		lon_0:long_name = "longitude" ;

// global attributes:
		:creation_date = "Mon Nov 13 22:47:49 MST 2017" ;
		:NCL_Version = "6.4.0" ;
		:system = "Linux geyser10 2.6.32-358.el6.x86_64 #1 SMP Wed Nov 2 11:00:18 MDT 2016 x86_64 x86_64 x86_64 GNU/Linux" ;
		:Conventions = "None" ;
		:grib_source = "gfs.0p25.2015012806.f000.grib2.tian267521.grb2" ;
		:title = "NCL: convert-GRIB-to-netCDF" ;
		:history = "Mon Nov 13 22:47:49 2017: ncks -O -d lat_0,3.0,54.0 -d lon_0,73.0,136.0 gfs.0p25.2015012806.f000.grib2.tian267521.nc gfs.0p25.2015012806.f000.grib2.tian267521.nc" ;
		:NCO = "4.4.2" ;
}
